    Mac OS X            	   2  �     �                                      ATTR      �  (   �                 (     com.apple.TextEncoding     7     com.apple.lastuseddate#PS      G   y  7com.apple.metadata:kMDLabel_voah4bcruwlmgbvk5fxagkek3q     �     com.apple.quarantine utf-8;134217984e3�h    ��O5    ��Ĭ�BG��[5��DΈ{D�#P�l�L����\�>�0�����6�T%����n��²�o@:��3��C|�)�o@h>�0f��^�T��y�ְ�� ���ح�|G�n!�t^�E4����q/0081;00000000;; 