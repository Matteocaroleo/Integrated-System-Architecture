    Mac OS X            	   2   �      �                                      ATTR       �   �                     �     com.apple.quarantine q/0081;6890d9ba;Telegram; 